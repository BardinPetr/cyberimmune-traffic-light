component trafficlight.CExternalControl

endpoints {
    ctrl : trafficlight.IExternalControl
    diag : trafficlight.IExternalDiagnostics
}