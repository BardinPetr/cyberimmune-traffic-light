component trafficlight.CTargetState

endpoints {
    stateInput : trafficlight.ITargetState
}