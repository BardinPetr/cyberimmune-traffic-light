component trafficlight.CExternalControl

endpoints {
    ctrl : trafficlight.IExternalControl
}