component trafficlight.CLightMode

endpoints {
    mode : trafficlight.ILightMode
}