component trafficlight.CDiagnostics

endpoints {
    diag : trafficlight.IDiagnostics
}